module main

// This file is just to help V recognize the project structure
// The actual framework code is in vwebx/server.v
fn main() {
    println('VWebX framework')
} 